-----------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Additional standard or custom libraries go here
entity comparator is
 generic(
 DATA_WIDTH : natural := 4
 );
port(
 --Inputs
 DINL : in std_logic_vector (DATA_WIDTH downto 0);
 DINR : in std_logic_vector (DATA_WIDTH - 1 downto 0);
 --Outputs
 DOUT : out std_logic_vector (DATA_WIDTH - 1 downto 0);
 isGreaterEq : out std_logic
 );
end entity comparator;
architecture behavioral of comparator is
--Signals and components go here
	signal intDINL : integer;
	signal intDINR : integer;
	
begin
	intDINL<=to_integer(unsigned(DINL));
	intDINR<=to_integer(unsigned(DINR));
	compute_diff: process(intDINL, intDINR)
		variable temp : integer;
	begin
		temp:=intDINL-intDINR;
		if (temp<0) then 
			DOUT<= DINL(DATA_WIDTH-1 downto 0);
			isGreaterEq<='0';
		else
			DOUT<=std_logic_vector(to_unsigned(temp,DATA_WIDTH));
			isGreaterEq<='1';
		end if;
	end process;
	
end architecture behavioral;

-----------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
--Additional standard or custom libraries go here
entity comparator is
 generic(
 DATA_WIDTH : natural := 4
 );
port(
 --Inputs
 DINL : in std_logic_vector (DATA_WIDTH downto 0);
 DINR : in std_logic_vector (DATA_WIDTH - 1 downto 0);
 --Outputs
 DOUT : out std_logic_vector (DATA_WIDTH - 1 downto 0);
 isGreaterEq : out std_logic
 );
end entity comparator;
architecture behavioral of comparator is
--Signals and components go here
begin
--Behavioral design goes here
end architecture behavioral;
----------------------------------------------------------------------------- 